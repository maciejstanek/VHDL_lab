library ieee;
use ieee.std_logic_1164.all;

entity counter_bcd_2digits is
  port(clk: in std_logic;
       digit_1: out std_logic_vector(6 downto 0);
       digit_10: out std_logic_vector(6 downto 0));
end entity counter_bcd_2digits;

architecture struct of counter_bcd_2digits is
begin
     
end architecture struct;    
