
* Project TESTING_SIGMA_DELTA
* Mentor Graphics Netlist Created with Version 5.10.3 Update-1
* File created Thu Apr 26 16:31:36 2018
* Inifile   : 
*
* Config file: C:\MentorGraphics\SystemVision5.10\standard\svspice.cfg
*
* Options   : -_ -h -kC:\MentorGraphics\SystemVision5.10\standard\svspice.cfg -gtesting_sigma_delta.tempfile 
* 
* Levels    : 
* 
.option noinclib
* Models for Eldo<->VHDL-AMS data conversion
.model a2d_eldo a2d mode=std_logic
.model d2a_eldo d2a mode=std_logic
.defhook a2d_eldo
.defhook d2a_eldo
YSUMMINGAMP5 SUMMINGAMP PORT: IN_A OUT2_A SUM2_A
YN1I107 ANALOG_INT(DEFAULT) PORT: SUM2_A N1N142
YN1I112 DAC_1B(DEFAULT) GENERIC: VMAX="-1.0" VMIN="1.0" PORT: OUT2_D OUT2_A
YN1I113 DECIM(DEFAULT) GENERIC: OSR="32" PORT: CLK OUT2_D DECIM2_A
YSUMMINGAMP6 SUMMINGAMP PORT: N1N142 OUT2_A N1N145
YN1I132 ANALOG_INT(DEFAULT) PORT: N1N145 N1N135
YN1I133 ADC_1B(DEFAULT) PORT: CLK N1N135 OUT2_D
YSUMMINGAMP4 SUMMINGAMP PORT: IN_A OUT_A SUM_A
YN1I72 ANALOG_INT(DEFAULT) PORT: SUM_A INT_SUM
YN1I75 ADC_1B(DEFAULT) PORT: CLK INT_SUM OUT_D
YN1I76 DAC_1B(DEFAULT) GENERIC: VMAX="-1.0" VMIN="1.0" PORT: OUT_D OUT_A
YCLOCK3 CLOCK(IDEAL) GENERIC: PERIOD="1 MS" PORT: CLK
YV_SINE3 V_SINE(IDEAL) GENERIC: AMPLITUDE="1.0" FREQ="2.0" PORT: IN_A 0
YN1I92 DECIM(DEFAULT) GENERIC: OSR="32" PORT: CLK OUT_D DECIM_A
* DICTIONARY 1
* GND = 0
*Note: Floating node DECIM2_A.
*Note: Floating node DECIM_A.
.GLOBAL ELECTRICAL_REF
.model DECIM(DEFAULT) macro lang=vhdlams LIB=WORK
.model SUMMINGAMP macro lang=vhdlams LIB=EDULIB
.model ANALOG_INT(DEFAULT) macro lang=vhdlams LIB=WORK
.model DAC_1B(DEFAULT) macro lang=vhdlams LIB=WORK
.model ADC_1B(DEFAULT) macro lang=vhdlams LIB=WORK
.model V_SINE(IDEAL) macro lang=vhdlams LIB=EDULIB
.model CLOCK(IDEAL) macro lang=vhdlams LIB=EDULIB
.END
